notes about FPGA 

A logic cell consists of a lookup table, a flip flop, and connection to adjacent cells. ... A logic slice consists of 2 logic cells. Xilinx counts closer to 2.25 logic cells per slice because they can do more per configurable logic block (CLB) than other architectures.

